`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////
// This file is a part of the Antarctic Impulsive Transient Antenna (ANITA)
// project, a collaborative scientific effort between multiple institutions. For
// more information, contact Peter Gorham (gorham@phys.hawaii.edu).
//
// All rights reserved.
//
// Author: Patrick Allison, Ohio State University (allison.122@osu.edu)
// Author:
// Author:
////////////////////////////////////////////////////////////////////////////////
module TOP_v38(
		input nADS,
		input WnR,
		input nRD,
		inout [31:0] LD,
		input [7:2] LA,
		input nCS2,
		input nCS3,
		output nREADY,
		output nBTERM,
		
		input BCLKO,
		output LCLK,
		input CLK125_P,
		input CLK125_N,
		input CMD_P,
		input CMD_N,
		input [3:0] HOLD_P,
		input [3:0] HOLD_N,
		input REF_P,
		input REF_N,
	
		input [7:0] A1TC,
		input [7:0] A2TC,
		input [7:0] A3TC,
		input [7:0] A4TC,
		input [7:0] VTRG_A1TC,
		input [7:0] VTRG_A2TC,
		input [7:0] VTRG_A3TC,
		input [7:0] VTRG_A4TC,
		
		output [7:0] L1_P,
		output [7:0] L1_N,
		
		// LAB innputs.
		output 		 A_GCK,
		output		 A_GCCLR,
		output		 A_RAMP,
		output [3:0] A_CS,
		output [7:0] A_S,
		output 		 A_SELMAIN,
		output 		 A_SELTAIL,
		output 		 A_NRUN,
		input 		 A_HITBUS,
		input 		 A_RCO,
		input [11:0] A_DAT,
		output		 A_TREF_P,
		output		 A_TREF_N,
		
		output 		 B_GCK,
		output		 B_GCCLR,
		output		 B_RAMP,
		output [3:0] B_CS,
		output [7:0] B_S,
		output 		 B_SELMAIN,
		output 		 B_SELTAIL,
		output 		 B_NRUN,
		input 		 B_HITBUS,
		input 		 B_RCO,
		input [11:0] B_DAT,
		output		 B_TREF_P,
		output		 B_TREF_N,

		output 		 C_GCK,
		output		 C_GCCLR,
		output		 C_RAMP,
		output [3:0] C_CS,
		output [7:0] C_S,
		output 		 C_SELMAIN,
		output 		 C_SELTAIL,
		output 		 C_NRUN,
		input 		 C_HITBUS,
		input 		 C_RCO,
		input [11:0] C_DAT,
		output		 C_TREF_P,
		output		 C_TREF_N,

		output 		 D_GCK,
		output		 D_GCCLR,
		output		 D_RAMP,
		output [3:0] D_CS,
		output [7:0] D_S,
		output 		 D_SELMAIN,
		output 		 D_SELTAIL,
		output 		 D_NRUN,
		input 		 D_HITBUS,
		input 		 D_RCO,
		input [11:0] D_DAT,
		output		 D_TREF_P,
		output		 D_TREF_N,
		
		output SCLK,
		output NSYNC,
		output [7:0] DIN,
		
		// Unuseds.
		output [3:0] CALSNH,
		output [3:0] TCS,
		output [3:0] RSS		
    );

	// Global clocks.
	
	wire clk33;
	wire clk100;
	wire clk125;
	wire clk250;
	wire clk250b;
	
	// Clock output.
	wire [3:0] TREF_P;
	wire [3:0] TREF_N;
	assign A_TREF_P = TREF_P[0]; assign A_TREF_N = TREF_N[0];
	assign B_TREF_P = TREF_P[1]; assign B_TREF_N = TREF_N[1];
	assign C_TREF_P = TREF_P[2]; assign C_TREF_N = TREF_N[2];
	assign D_TREF_P = TREF_P[3]; assign D_TREF_N = TREF_N[3];
	
	// Reference pulse from TURF.
	wire REF;
	
	// TURF HOLD inputs
	wire [3:0] HOLD;

	// Global reset.
	
	wire clr_all;

	// MESSv2 <-> LAB_TOPv2 interface.
	wire [3:0] 		lab_digitize;
	wire [12:0] 	lab_addr;
	wire [31:0] 	lab_dat;
	wire 				lab_ready;

	// Trigger inputs.
	// These are NOT individual antennas. They're individual SHORT inputs.
	// At some point in the long, distant past, they were individual antennas.
	wire [7:0] ANT_A;
	wire [7:0] ANT_B;
	wire [7:0] ANT_C;
	wire [7:0] ANT_D;
	wire [31:0] trig_scaler_path;

	// Trigger outputs.
	wire [3:0] L1;
	// Uh... stuff, I guess.
	wire [31:0] CR;
	// Mask register, I guess?
	wire [31:0] short_mask;
	// Some monitoring stuff that I have no idea what it does.
	wire [7:0] mon_scaler;
	wire L1MON2;
	wire L1MON3;
	wire L1MON4;
	
	SURF_infrastructure #(.REF_CLOCK("125MHZ")) u_infrastructure( .clk33_o(clk33),
																					 .clk100_o(clk100),
																					 .clk125_o(clk125),
																					 .clk250_o(clk250),
																					 .clk250b_o(clk250b),
																					 .clr_all_i(clr_all),
																					 .CLK125_P(CLK125_P),.CLK125_N(CLK125_N),
																					 .LCLK(LCLK),
																					 .BCLKO(BCLKO),
																					 .CMD_P(CMD_P),.CMD_N(CMD_N),.CMD(command),
																					 .HOLD_P(HOLD_P),.HOLD_N(HOLD_N),.HOLD(HOLD),
																					 .TREF_P(TREF_P),.TREF_N(TREF_N),
																					 .REF_P(REF_P),.REF_N(REF_N),.REF(REF),
																					 .L1_P(L1_P),.L1_N(L1_N),.L1(L1));
	// Trigger infrastructure.
	Trig_RX u_trigger_rx(.A1TC(A1TC),.A2TC(A2TC),.A3TC(A3TC),.A4TC(A4TC),
								.VTRG_A1TC(VTRG_A1TC),.VTRG_A2TC(VTRG_A2TC),.VTRG_A3TC(VTRG_A3TC),.VTRG_A4TC(VTRG_A4TC),
								.out_for_scaler(trig_scaler_path),
								.ANT_A(ANT_A),.ANT_B(ANT_B),.ANT_C(ANT_C),.ANT_D(ANT_D));
	// Trigger.
	Level1_Trigger level1trigger(.ANT_A(ANT_A),.ANT_B(ANT_B),.ANT_C(ANT_C),.ANT_D(ANT_D),
									 .ANT_A_for_scalers(trig_scaler_path[0 +: 8]),
									 .ANT_B_for_scalers(trig_scaler_path[8 +: 8]),
									 .ANT_C_for_scalers(trig_scaler_path[16 +: 8]),
									 .ANT_D_for_scalers(trig_scaler_path[24 +: 8]),
									 .CLK(clk33),.CLR_ALL(clr_all),.REFPULSE(REF),								 
									 .L1(L1),
									 .mask_pass(short_mask),
									 .CR(CR),
									 .MONSCALER(mon_scaler),
									 .MON2(L1MON2),
									 .MON3(L1MON3),
									 .MON4(L1MON4),
									 .CLK125(clk125),
									 .CLK250(clk250),
									 .CLK250_180(clk250b));									 

	reg mon_bit = 0;
	reg mon_bit_clk33 = 0;
	reg mon_bit_clear = 0;
	always @(posedge clk250) begin
		if (CR[8]) mon_bit <= 1;
		else if (mon_bit_clear) mon_bit <= 0;
	end
	always @(posedge clk33) begin
		mon_bit_clk33 <= mon_bit;
		mon_bit_clear <= mon_bit_clk33;
	end
	
	wire [34:0] lab_debug;

	// LAB readout and memory.
	LAB_TOPv2 u_labtop( .clk_i(clk33),
							  .clk100_i(clk100),
							  .rst_i(clr_all),
							  .hold_i(HOLD),
							  .digitize_i(lab_digitize),
							  .addr_i(lab_addr),
							  .dat_o(lab_dat),
							  .done_o(lab_ready),
							  .A_SELTAIL(A_SELTAIL),
							  .A_SELMAIN(A_SELMAIN),
							  .A_GCK(A_GCK),
							  .A_RAMP(A_RAMP),
							  .A_GCCLR(A_GCCLR),
							  .A_NRUN(A_NRUN),
							  .A_CS(A_CS),
							  .A_S(A_S),
							  .A_HITBUS(A_HITBUS),
							  .A_RCO(A_RCO),
							  .A_DAT(A_DAT),
							  
							  .B_SELTAIL(B_SELTAIL),
							  .B_SELMAIN(B_SELMAIN),
							  .B_GCK(B_GCK),
							  .B_RAMP(B_RAMP),
							  .B_GCCLR(B_GCCLR),
							  .B_NRUN(B_NRUN),
							  .B_CS(B_CS),
							  .B_S(B_S),
							  .B_HITBUS(B_HITBUS),
							  .B_RCO(B_RCO),
							  .B_DAT(B_DAT),

							  .C_SELTAIL(C_SELTAIL),
							  .C_SELMAIN(C_SELMAIN),
							  .C_GCK(C_GCK),
							  .C_RAMP(C_RAMP),
							  .C_GCCLR(C_GCCLR),
							  .C_NRUN(C_NRUN),
							  .C_CS(C_CS),
							  .C_S(C_S),
							  .C_HITBUS(C_HITBUS),
							  .C_RCO(C_RCO),
							  .C_DAT(C_DAT),

							  .D_SELTAIL(D_SELTAIL),
							  .D_SELMAIN(D_SELMAIN),
							  .D_GCK(D_GCK),
							  .D_RAMP(D_RAMP),
							  .D_GCCLR(D_GCCLR),
							  .D_NRUN(D_NRUN),
							  .D_CS(D_CS),
							  .D_S(D_S),
							  .D_HITBUS(D_HITBUS),
							  .D_RCO(D_RCO),
							  .D_DAT(D_DAT),
							  .debug_o(lab_debug)
		);


	wire dac_wr;
	wire dac_busy;
	wire dac_update;
	wire [4:0] dac_waddr;
	wire [4:0] dac_raddr;
	wire [15:0] dac_dat_in;
	wire [15:0] dac_dat_out;

	wire [34:0] td_debug;
	assign td_debug[0] = mon_bit_clear;
	assign td_debug[1 +: 8] = DIN;
	assign td_debug[9] = SCLK;
	assign td_debug[10] = NSYNC;
	assign td_debug[11] = dac_wr;
	assign td_debug[12 +: 12] = dac_dat_in;
	assign td_debug[24 +: 4] = dac_waddr;
	assign td_debug[28] = dac_update;
	assign td_debug[29] = dac_busy;

	DAC_CTRL_v3 u_dacs( 	.clk_i(clk33),
								.dac_we_i(dac_wr),
								.busy_o(dac_busy),
								.dac_waddr_i(dac_waddr),
								.dac_dat_i(dac_dat_in),
								.dac_raddr_i(dac_raddr),
								.dac_dat_o(dac_dat_out),
								.update_i(dac_update),
								.SCLK(SCLK),
								.NSYNC(NSYNC),
								.DIN(DIN));
								

	// MESS debugging.
	wire [34:0] debug;
	wire [4:0] rfp_addr;
	// PLX/register interface
	MESSv2 u_mess(		  .clk_i(clk33),
							  .cmd_i(command),
							  .lab_dat_i(lab_dat),
							  .lab_ready_i(lab_ready),
							  .lab_addr_o(lab_addr),
							  .lab_digitize_o(lab_digitize),

							  .rfp_dat_i(rfp_addr),
							  .rfp_addr_o(rfp_addr),
							  .clr_all_o(clr_all),

							  .dac_waddr_o(dac_waddr),
							  .dac_raddr_o(dac_raddr),
							  .dac_wr_o(dac_wr),
							  .dac_update_o(dac_update),
							  .dac_busy_i(dac_busy),
							  .dac_dat_i(dac_dat_out),
							  .dac_dat_o(dac_dat_in),
							  
							  .short_mask_o(short_mask),
							  
							  .nADS(nADS),
							  .WnR(WnR),
							  .LA(LA),
							  .LD(LD),
							  .nCS2(nCS2),
							  .nCS3(nCS3),
							  .nRD(nRD),
							  .nREADY(nREADY),
							  .nBTERM(nBTERM),
							  .debug_o(debug)
	);
	
	// ChipScope debugging cores.
	wire [35:0] ila_control;
	(* BOX_TYPE = "black_box" *)
	cs_icon u_icon(.CONTROL0(ila_control));
	(* BOX_TYPE = "black_box" *)
	cs_ila u_ila(.CONTROL(ila_control),.CLK(clk33),.TRIG0(debug));

	// Unused LAB test crap.
	// CALSNH = VCC
	// RSS = VCC
	// TCS = GND
	assign CALSNH = {4{1'b1}};
	assign RSS = {4{1'b1}};
	assign TCS = {4{1'b0}};
	
endmodule
